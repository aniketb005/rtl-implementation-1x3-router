/************************************************************************

 Copyright 2019 - Maven Silicon Softech Pvt Ltd.  
 
 www.maven-silicon.com
 
 All Rights Reserved
   
 This source code is an unpublished work belongs to Maven Silicon Softech Pvt Ltd.
 It is not to be shared with or used by any third parties who have not enrolled for our
 paid training courses or received any written authorization from Maven Silicon.

Filename:	ram_test_pkg.sv   

Version:	1.0

************************************************************************/
package test_pkg;


//import uvm_pkg.sv
	import uvm_pkg::*;
//include uvm_macros.sv
	`include "uvm_macros.svh"
`include "tb_defs.sv"
`include "write_xtn.sv"
`include "wr_agent_config.sv"
`include "rd_agent_config.sv"
`include "env_config.sv"
`include "wr_driver.sv"
`include "wr_monitor.sv"
`include "wr_sequencer.sv"
`include "wr_agent.sv"
`include "wr_agt_top.sv"
`include "wr_seqs.sv"

`include "read_xtn.sv"
`include "rd_monitor.sv"
`include "rd_sequencer.sv"
`include "rd_seqs.sv"
`include "rd_driver.sv"
`include "rd_agent.sv"
`include "rd_agt_top.sv"

`include "virtual_sequencer.sv"
`include "virtual_seqs.sv"
`include "scoreboard.sv"

`include "tb.sv"


`include "vtest_lib.sv"
endpackage
